library verilog;
use verilog.vl_types.all;
entity PIPELINE_IF_ID_vlg_vec_tst is
end PIPELINE_IF_ID_vlg_vec_tst;
