library verilog;
use verilog.vl_types.all;
entity Data_memory_diagram_vlg_check_tst is
    port(
        Read_data       : in     vl_logic_vector(7 downto 0);
        sampler_rx      : in     vl_logic
    );
end Data_memory_diagram_vlg_check_tst;
