library verilog;
use verilog.vl_types.all;
entity Processor_MIPS_with_Pipelines_diagram_vlg_vec_tst is
end Processor_MIPS_with_Pipelines_diagram_vlg_vec_tst;
