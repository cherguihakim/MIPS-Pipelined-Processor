library verilog;
use verilog.vl_types.all;
entity DECODEUR_3_x_8_vlg_check_tst is
    port(
        sortie_0        : in     vl_logic;
        sortie_1        : in     vl_logic;
        sortie_2        : in     vl_logic;
        sortie_3        : in     vl_logic;
        sortie_4        : in     vl_logic;
        sortie_5        : in     vl_logic;
        sortie_6        : in     vl_logic;
        sortie_7        : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end DECODEUR_3_x_8_vlg_check_tst;
