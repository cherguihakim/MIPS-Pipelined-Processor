library verilog;
use verilog.vl_types.all;
entity TEST_CONTROL_ALU_vlg_vec_tst is
end TEST_CONTROL_ALU_vlg_vec_tst;
