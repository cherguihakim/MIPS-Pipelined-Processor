library verilog;
use verilog.vl_types.all;
entity Instruction_memory_diagram_vlg_vec_tst is
end Instruction_memory_diagram_vlg_vec_tst;
