library verilog;
use verilog.vl_types.all;
entity CONTROL_PC_vlg_check_tst is
    port(
        selecteur_PC    : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end CONTROL_PC_vlg_check_tst;
