library verilog;
use verilog.vl_types.all;
entity FORWARDING_UNIT_vlg_vec_tst is
end FORWARDING_UNIT_vlg_vec_tst;
