library verilog;
use verilog.vl_types.all;
entity DECODEUR_3_x_8_vlg_vec_tst is
end DECODEUR_3_x_8_vlg_vec_tst;
