INSTRUCTION_MEMORY_inst : INSTRUCTION_MEMORY PORT MAP (
		address	 => address_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
