LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ALU_CONTROL IS 
PORT(ALU_OP : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
     FUNCTION_CODE : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
     SEL_ALU : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)   );
END ALU_CONTROL;

ARCHITECTURE STRUCT OF ALU_CONTROL IS 

BEGIN

SEL_ALU(2) <= (ALU_OP(0)) OR (ALU_OP(1) AND FUNCTION_CODE(1));

SEL_ALU(1) <= (NOT(ALU_OP(1))) OR NOT((FUNCTION_CODE(2)));

SEL_ALU(0) <= (ALU_OP(1)) AND (FUNCTION_CODE(3) OR FUNCTION_CODE(0));

END STRUCT;