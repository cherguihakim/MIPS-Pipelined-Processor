library verilog;
use verilog.vl_types.all;
entity REGISTER_FILE_vlg_vec_tst is
end REGISTER_FILE_vlg_vec_tst;
