library verilog;
use verilog.vl_types.all;
entity ALU_8BITS_vlg_vec_tst is
end ALU_8BITS_vlg_vec_tst;
