library verilog;
use verilog.vl_types.all;
entity BIG_MUX_vlg_vec_tst is
end BIG_MUX_vlg_vec_tst;
