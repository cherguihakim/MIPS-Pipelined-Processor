library verilog;
use verilog.vl_types.all;
entity Diagram_test_sans_PC_vlg_vec_tst is
end Diagram_test_sans_PC_vlg_vec_tst;
