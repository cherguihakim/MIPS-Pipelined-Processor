library verilog;
use verilog.vl_types.all;
entity HAZARD_UNIT_vlg_vec_tst is
end HAZARD_UNIT_vlg_vec_tst;
