library verilog;
use verilog.vl_types.all;
entity five_bit_comparator_vlg_vec_tst is
end five_bit_comparator_vlg_vec_tst;
