library verilog;
use verilog.vl_types.all;
entity CONTROL_PC_vlg_vec_tst is
end CONTROL_PC_vlg_vec_tst;
