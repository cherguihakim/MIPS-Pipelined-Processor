library verilog;
use verilog.vl_types.all;
entity register8bits_affichage_vlg_vec_tst is
end register8bits_affichage_vlg_vec_tst;
